LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY main IS
 GENERIC(W : NATURAL := 18);
 PORT (
 IS_ON : IN BIT; -- Indica se est� ligado.
 MODE : IN BIT; -- Aumenta ou n�o o slp
 UP : IN BIT; -- Incrementa o contador atual
 DOWN : IN BIT; -- Decrementa o contador atual
 SLEEP : IN BIT; -- Bot�o de soneca
 CLK : IN BIT; -- Clock
 HorasDezenas : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
 HorasUnidades : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
 MinutosDezenas : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
 MinutosUnidades : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
 );
END main;

-----------------------------------------------------------

ARCHITECTURE Behavior OF main IS

COMPONENT demux_2x1 IS
GENERIC (W : NATURAL := 18);
PORT (
  s : IN BIT;
  sel : IN BIT;
  a, b : OUT BIT
);
END COMPONENT;

COMPONENT mux_2x1 IS
GENERIC (W : NATURAL := 18);
PORT (a, b : IN BIT_VECTOR (W-1 DOWNTO 0);
       sel : IN BIT;
         s : OUT BIT_VECTOR (W-1 DOWNTO 0));
END COMPONENT;

COMPONENT comparador IS
   GENERIC (W : NATURAL := 18);
   PORT (e1, e2: IN STD_LOGIC_VECTOR (W-1 DOWNTO 0);
         saida : OUT STD_LOGIC);
END COMPONENT;

COMPONENT counter_18bits IS
 GENERIC(W : NATURAL := 18);
 PORT (
   clk : IN BIT; -- clock
   clrn: IN BIT; -- clear
   ena : IN BIT; -- enable
   q : BUFFER STD_LOGIC_VECTOR(W-1 DOWNTO 0)
 );
END COMPONENT;

COMPONENT Divider is
GENERIC(W : NATURAL := 18);
port(
  X   : in STD_LOGIC_VECTOR(W-1 downto 0);
  Y   : in STD_LOGIC_VECTOR(W-1 downto 0);
  R   : out STD_LOGIC_VECTOR(W-1 downto 0)
);
END COMPONENT;

COMPONENT offset_mem IS
 GENERIC(W : NATURAL := 18);
 PORT (
   is_on : IN BIT;
   up : IN BIT;
   down: IN BIT;
   q : BUFFER STD_LOGIC_VECTOR(W-1 DOWNTO 0)
 );
END COMPONENT;

COMPONENT sleep_offset IS
 GENERIC(W : NATURAL := 18);
 PORT (
 increase : IN BIT; -- aumenta ou n�o o slp
 reset : IN BIT; -- reseta o slp
 q : BUFFER STD_LOGIC_VECTOR(W-1 DOWNTO 0));
END COMPONENT;

COMPONENT alarm_counter IS
 GENERIC(W : NATURAL := 18);
 PORT (
 start : IN BIT; -- clear
 kill : BUFFER BIT; -- clock
 q : BUFFER STD_LOGIC_VECTOR(W-1 DOWNTO 0));
END COMPONENT;

COMPONENT encoder_bin_to_dec IS
PORT( din : IN STD_LOGIC_VECTOR(17 DOWNTO 0); -- DATA IN
      dout : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) ); -- DATA OUT
END COMPONENT;

COMPONENT decoder_dec_to_display IS
PORT( din : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- DATA INPUT
      display : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT;

------------------------------------------------------------
-- SIGNAL IS_OFF : BIT;
SIGNAL TOTALMAXSECONDS : STD_LOGIC_VECTOR(W-1 DOWNTO 0);

SIGNAL CLOCK1OUT : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL CLOCK2OUT : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL TEMPCLOCKTIME : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL CLOCKTIME : STD_LOGIC_VECTOR(W-1 DOWNTO 0);

SIGNAL ALARMOUT1 : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL ALARMOUT2 : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL TEMPALARMTIME : STD_LOGIC_VECTOR(W-1 DOWNTO 0);
SIGNAL ALARMTIME : STD_LOGIC_VECTOR(W-1 DOWNTO 0);

SIGNAL TODISPLAY : STD_LOGIC_VECTOR(W-1 DOWNTO 0);

SIGNAL CLOCKUP : BIT;
SIGNAL CLOCKDOWN : BIT;
SIGNAL ALARMUP : BIT;
SIGNAL ALARMDOWN : BIT;

SIGNAL ALARM_COUNT_IS_OVER : BIT;
SIGNAL ALARM_FLAG : BIT;

BEGIN
  
  TOTALMAXSECONDS <= "010101000110000000";
  
  updemux : demux_2x1
    PORT MAP( UP, MODE, CLOCKUP, ALARMUP );
      
  downdemux : demux_2x1
    PORT MAP( DOWN, MODE, CLOCKDOWN, ALARMDOWN );
      
  clock1 : counter_18bits
    PORT MAP( CLK, IS_ON, IS_ON, CLOCK1OUT );

  clock2 : offset_mem
    PORT MAP( IS_ON, CLOCKUP, CLOCKDOWN, CLOCK2OUT );
      
  alarm1 : offset_mem
    PORT MAP( IS_ON, ALARMUP, ALARMDOWN, ALARMOUT1 );
  
  alarmcnt : alarm_counter
    PORT MAP( CLK, [strt], [KIL], [ALARMOUT2] );
  
  alarm2 : sleep_offser
    PORT MAP([KIL_OLD], ![NOT_EMPTY], ALARMOUT2 );
      
  TEMPCLOCKTIME <= CLOCKOUT1 + CLOCKOUT2;
  CLOCKTIME <= STD_LOGIC_VECTOR( unsigned(TEMPCLOCKTIME) mod unsigned(TOTALMAXSECONDS) );
  
  TEMPALARMTIME <= ALARMOUT1 + ALARMOUT2;
  ALARMTIME <= STD_LOGIC_VECTOR( unsigned(TEMPALARMTIME) mod unsigned(TOTALMAXSECONDS) );
      
  ALARM_COUNT_IS_OVER <= ( ALARMOUT2 = "000000000000000000" );
  
  ALARM_FLAG <= ( CLOCKTIME = ALARMTIME );
  
  display_mux : mux_2x1
    PORT MAP( CLOCKTIME, ALARMTIME, MODE, TODISPLAY );
  
  
      
  
      
END Behavior;
